library IEEE;
use IEEE.std_logic_1164.all;

entity and is
    port(
        a, b: in std_logic;
        c   : out std_logic
    );
end and;

architecture behave of and is
begin
    c <= a and b;
end behave;